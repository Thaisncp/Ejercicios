library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity ejercicio22 is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           S1 : out  STD_LOGIC;
           S2 : out  STD_LOGIC;
           S3 : out  STD_LOGIC);
end ejercicio22;

architecture sensor of ejercicio22 is

begin
	S1 <= '1' when (A = '0' and B = '0');
	S2 <= '1' when (A = '1' and B = '1');
	S3 <= '1' when (A = '1' and B = '1');
end sensor;
