library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity entidad2 is
    Port ( A : in  STD_LOGIC;
           B : in  STD_LOGIC;
           C : out  STD_LOGIC);
end entidad2;

