library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity vectores2 is
	port (A : in std_logic_vector(0 to 3);
	 	B : in std_logic_vector(0 to 3);
		C : out std_logic_vector(0 to 3));
end vectores2;


