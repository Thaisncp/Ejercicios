library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity circuito2 is
	port(a : in bit_vector(0 to 3)
		   b : in bit_vector(0 to 3)
		   f : out std_logic);
end circuito2;
