library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity entidad is
    Port ( P0 : in  STD_LOGIC;
           P1 : in  STD_LOGIC;
           P2 : in  STD_LOGIC;
           A0 : out  STD_LOGIC;
           A1 : out  STD_LOGIC;
           X : inout  STD_LOGIC);
end entidad;
